module background( input                             Clk,
                    output logic [0:11][0:143][0:5]  dive_health_bar, kick_health_bar,
					output logic [0:19][0:199][0:5]     p1_win, p2_win,
                    output logic [0:39][0:199][0:5]     title
				 );

    always_comb
    begin
        dive_health_bar <=
        '{
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,61,0,0,0,0,0,61,61,0,0,61,61,0,0,0,0,61,61,0,0,61,61,61,61,61,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,61,61,61,0,0,0,61,61,0,0,61,61,0,0,0,0,61,61,0,0,61,61,61,61,61,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,0,61,61,61,0,0,61,61,0,0,0,61,61,0,0,61,61,0,0,0,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,0,0,61,61,0,0,61,61,0,0,0,61,61,0,0,61,61,0,0,0,61,61,61,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,0,0,61,61,0,0,61,61,0,0,0,0,61,61,61,61,0,0,0,0,61,61,61,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,0,61,61,61,0,0,61,61,0,0,0,0,61,61,61,61,0,0,0,0,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,61,61,61,0,0,0,61,61,0,0,0,0,0,61,61,0,0,0,0,0,61,61,61,61,61,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,61,61,61,0,0,0,0,0,61,61,0,0,0,0,0,61,61,0,0,0,0,0,61,61,61,61,61,61,61,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
        };

        kick_health_bar <=
        '{
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,0,0,61,0,0,61,61,61,61,61,61,0,0,0,0,61,61,0,0,61,61,0,0,61,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,0,61,61,0,0,61,61,61,61,61,61,0,0,61,61,61,61,0,0,61,61,0,61,61,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,61,61,0,0,0,0,0,61,61,0,0,0,0,61,61,0,0,0,0,61,61,61,61,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,61,0,0,0,0,0,0,61,61,0,0,0,0,61,61,0,0,0,0,61,61,61,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,61,61,0,0,0,0,0,61,61,0,0,0,0,61,61,0,0,0,0,61,61,61,61,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,61,61,0,0,0,0,0,61,61,0,0,0,0,61,61,0,0,0,0,61,61,61,61,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,0,61,61,0,0,61,61,61,61,61,61,0,0,61,61,61,61,0,0,61,61,0,61,61,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,61,61,0,61,61,0,0,61,61,61,61,61,61,0,0,0,0,61,61,0,0,61,61,0,61,61,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
        };

        p1_win <=
'{
'{55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,55,55,56,56,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,56,56,56,56,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55,56,56,56,56,55,55,55,55,55,55,56,56,56,56,55,55,56,56,56,56,55,55,56,56,56,56,55,55,55,55,56,56,56,56,55,55,55,55,56,56,56,56,56,56,56,56,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55}
};

        p2_win <=
'{
'{55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,55,55,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,57,57,55,55,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,57,57,55,55,57,57,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,57,57,55,55,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,57,57,57,57,57,57,55,55,57,57,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,57,57,57,57,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55,55,55,57,57,57,57,55,55,55,55,55,55,57,57,57,57,55,55,57,57,57,57,55,55,57,57,57,57,55,55,55,55,57,57,57,57,55,55,55,55,57,57,57,57,57,57,57,57,55,55,55,55,55,55,55,55},
'{55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55}
};

        title <=
'{
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,0,0,0,0,0,0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0,0,0,54,54,54,54,54,54,54,54,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};

    end
endmodule